----------------------------------------------------------------------------------
-- Engineer: pedram babakhani
-- 
-- Create Date: 09/04/2017 06:19:37 PM
-- Design Name: 
-- Module Name: LSTM_TB - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


LIBRARY IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.ALL;
LIBRARY WORK;
USE IEEE.std_logic_textio.all;
USE WORK.Generic_size_of_matrices_pkg.ALL;
library std;
use std.textio.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

ENTITY LSTM_TB is
--  Port ( );
END LSTM_TB;

ARCHITECTURE Behavioral OF LSTM_TB IS


SIGNAL CLK_tb : STD_LOGIC :='0';
SIGNAL RST_tb : STD_LOGIC;  
SIGNAL EN_tb : STD_LOGIC;   
SIGNAL Done_tb : STD_LOGIC;                
SIGNAL X_t_tb :  Fixed_Point; -- X(t)
SIGNAL H_t1_tb : Fixed_Point; -- H(t-1)
SIGNAL C_t1_tb : Fixed_Point; -- C(t-1)
SIGNAL H_t_tb :  Fixed_Point; -- H(t)
SIGNAL C_t_tb :  Fixed_Point; -- C(t)
CONSTANT half_period : Time:= 5ns;
CONSTANT period : Time:= 10ns;
SIGNAL flag : STD_LOGIC := '0';  

COMPONENT LSTM_Core  
            PORT ( 
            CLK : IN STD_LOGIC; -- Clock
            RST : IN STD_LOGIC; -- Reset
            En : IN STD_LOGIC; -- Enable
            X_t : IN Fixed_Point; -- X(t)
            H_t1 : IN Fixed_Point; -- H(t-1)
            C_t1 : IN Fixed_Point; -- C(t-1)
            H_t : OUT Fixed_Point; -- H(t)
            C_t : OUT Fixed_Point; -- C(t)
            Done : OUT STD_LOGIC); --Done
END COMPONENT;
 
BEGIN
DUT : LSTM_Core
  PORT MAP (
    CLK => CLK_tb,
    RST => RST_tb,
    EN => En_tb,
    X_t =>   X_t_tb,
    H_t1 => H_t1_tb,
    C_t1 => C_t1_tb,
    H_t =>   H_t_tb,
    C_t =>   C_t_tb,
    Done => Done_tb);
    

 CLK_tb <= NOT CLK_tb AFTER half_period;   
 
 X_t_tb <=  ("00000000000000010000000000000000"), 
 ("00000000000000000000000000000000") AFTER 10ns, 
 ("00000000000000010000000000000000") AFTER 20ns,
 ("00000000000000000000000000000000") AFTER 30ns,
 ("00000000000000000000000000000000") AFTER 40ns,
 ("00000000000000000000000000000000") AFTER 50ns,
 ("00000000000000010000000000000000") AFTER 60ns,
 ("00000000000000000000000000000000") AFTER 70ns,
 ("00000000000000000000000000000000") AFTER 80ns,
 ("00000000000000000000000000000000") AFTER 90ns,
 ("00000000000000010000000000000000") AFTER 10ns,
 ("00000000000000000000000000000000") AFTER 110ns,
 ("00000000000000000010000111001100") AFTER 120ns,
 ("00000000000000000000000000000000") AFTER 130ns,
 ("00000000000000000000000000000000") AFTER 140ns,
 ("00000000000000000000000000000000") AFTER 150ns,
 ("00000000000000000000000000000000") AFTER 160ns,
 ("00000000000000000000000000000000") AFTER 170ns,
 ("00000000000000010000000000000000") AFTER 180ns,
 ("00000000000000010000000000000000") AFTER 190ns,
 ("00000000000000010000000000000000") AFTER 200ns,
 ("00000000000000000000000000000000") AFTER 210ns,
 ("00000000000000000000000000000000") AFTER 220ns,
 ("00000000000000000000000000000000") AFTER 230ns,
 ("00000000000000010000000000000000") AFTER 240ns,
 ("00000000000000000000000000000000") AFTER 250ns,
 ("00000000000000010000000000000000") AFTER 260ns;

 H_t1_tb <=  ("00000000000000000000000000000000"),
 ("00000000000000000000000000000000")  AFTER 10ns,   
 ("00000000000000000000000000000000")  AFTER 20ns,   
 ("00000000000000000000000000000000")  AFTER 30ns,   
 ("00000000000000000000000000000000")  AFTER 40ns,   
 ("00000000000000000000000000000000")  AFTER 50ns,   
 ("00000000000000000000000000000000")  AFTER 60ns,   
 ("00000000000000000000000000000000")  AFTER 70ns,   
 ("00000000000000000000000000000000")  AFTER 80ns,   
 ("00000000000000000000000000000000")  AFTER 90ns,   
 ("00000000000000000000000000000000")  AFTER 10ns,   
 ("00000000000000000000000000000000")  AFTER 110ns,  
 ("00000000000000000000000000000000")  AFTER 120ns,  
 ("00000000000000000000000000000000")  AFTER 130ns,  
 ("00000000000000000000000000000000")  AFTER 140ns,  
 ("00000000000000000000000000000000")  AFTER 150ns,  
 ("00000000000000000000000000000000")  AFTER 160ns,  
 ("00000000000000000000000000000000")  AFTER 170ns,  
 ("00000000000000000000000000000000")  AFTER 180ns,  
 ("00000000000000000000000000000000")  AFTER 190ns,  
 ("00000000000000000000000000000000")  AFTER 200ns,  
 ("00000000000000000000000000000000")  AFTER 210ns,  
 ("00000000000000000000000000000000")  AFTER 220ns,  
 ("00000000000000000000000000000000")  AFTER 230ns,  
 ("00000000000000000000000000000000")  AFTER 240ns,  
 ("00000000000000000000000000000000")  AFTER 250ns,  
 ("00000000000000000000000000000000")  AFTER 260ns,  
 ("00000000000000000000000000000000")  AFTER 270ns,  
 ("00000000000000000000000000000000")  AFTER 280ns,  
 ("00000000000000000000000000000000")  AFTER 290ns,  
 ("00000000000000000000000000000000")  AFTER 300ns,  
 ("00000000000000000000000000000000")  AFTER 310ns,  
 ("00000000000000000000000000000000")  AFTER 320ns,  
 ("00000000000000000000000000000000")  AFTER 330ns,  
 ("00000000000000000000000000000000")  AFTER 340ns,  
 ("00000000000000000000000000000000")  AFTER 350ns,  
 ("00000000000000000000000000000000")  AFTER 360ns,  
 ("00000000000000000000000000000000")  AFTER 370ns,  
 ("00000000000000000000000000000000")  AFTER 380ns,  
 ("00000000000000000000000000000000")  AFTER 390ns,  
 ("00000000000000000000000000000000")  AFTER 400ns,  
 ("00000000000000000000000000000000")  AFTER 410ns,  
 ("00000000000000000000000000000000")  AFTER 420ns,  
 ("00000000000000000000000000000000")  AFTER 430ns,  
 ("00000000000000000000000000000000")  AFTER 440ns,  
 ("00000000000000000000000000000000")  AFTER 450ns,  
 ("00000000000000000000000000000000")  AFTER 460ns,  
 ("00000000000000000000000000000000")  AFTER 470ns,  
 ("00000000000000000000000000000000")  AFTER 480ns,  
 ("00000000000000000000000000000000")  AFTER 490ns,  
 ("00000000000000000000000000000000")  AFTER 500ns,  
 ("00000000000000000000000000000000")  AFTER 510ns,  
 ("00000000000000000000000000000000")  AFTER 520ns,  
 ("00000000000000000000000000000000")  AFTER 530ns,  
 ("00000000000000000000000000000000")  AFTER 540ns,
 ("00000000000000000000000000000000")  AFTER 550ns;  


 C_t1_tb <=  ("00000000000000000000000000000000"),
 ("00000000000000000000000000000000") AFTER 10ns,  
 ("00000000000000000000000000000000") AFTER 20ns,  
 ("00000000000000000000000000000000") AFTER 30ns,  
 ("00000000000000000000000000000000") AFTER 40ns,  
 ("00000000000000000000000000000000") AFTER 50ns,  
 ("00000000000000000000000000000000") AFTER 60ns,  
 ("00000000000000000000000000000000") AFTER 70ns,  
 ("00000000000000000000000000000000") AFTER 80ns,  
 ("00000000000000000000000000000000") AFTER 90ns,  
 ("00000000000000000000000000000000") AFTER 10ns,  
 ("00000000000000000000000000000000") AFTER 110ns, 
 ("00000000000000000000000000000000") AFTER 120ns, 
 ("00000000000000000000000000000000") AFTER 130ns, 
 ("00000000000000000000000000000000") AFTER 140ns, 
 ("00000000000000000000000000000000") AFTER 150ns, 
 ("00000000000000000000000000000000") AFTER 160ns, 
 ("00000000000000000000000000000000") AFTER 170ns, 
 ("00000000000000000000000000000000") AFTER 180ns, 
 ("00000000000000000000000000000000") AFTER 190ns, 
 ("00000000000000000000000000000000") AFTER 200ns, 
 ("00000000000000000000000000000000") AFTER 210ns, 
 ("00000000000000000000000000000000") AFTER 220ns, 
 ("00000000000000000000000000000000") AFTER 230ns, 
 ("00000000000000000000000000000000") AFTER 240ns, 
 ("00000000000000000000000000000000") AFTER 250ns, 
 ("00000000000000000000000000000000") AFTER 260ns, 
 ("00000000000000000000000000000000") AFTER 270ns, 
 ("00000000000000000000000000000000") AFTER 280ns, 
 ("00000000000000000000000000000000") AFTER 290ns, 
 ("00000000000000000000000000000000") AFTER 300ns, 
 ("00000000000000000000000000000000") AFTER 310ns, 
 ("00000000000000000000000000000000") AFTER 320ns, 
 ("00000000000000000000000000000000") AFTER 330ns, 
 ("00000000000000000000000000000000") AFTER 340ns, 
 ("00000000000000000000000000000000") AFTER 350ns, 
 ("00000000000000000000000000000000") AFTER 360ns, 
 ("00000000000000000000000000000000") AFTER 370ns, 
 ("00000000000000000000000000000000") AFTER 380ns, 
 ("00000000000000000000000000000000") AFTER 390ns, 
 ("00000000000000000000000000000000") AFTER 400ns, 
 ("00000000000000000000000000000000") AFTER 410ns, 
 ("00000000000000000000000000000000") AFTER 420ns, 
 ("00000000000000000000000000000000") AFTER 430ns, 
 ("00000000000000000000000000000000") AFTER 440ns, 
 ("00000000000000000000000000000000") AFTER 450ns, 
 ("00000000000000000000000000000000") AFTER 460ns, 
 ("00000000000000000000000000000000") AFTER 470ns, 
 ("00000000000000000000000000000000") AFTER 480ns, 
 ("00000000000000000000000000000000") AFTER 490ns, 
 ("00000000000000000000000000000000") AFTER 500ns, 
 ("00000000000000000000000000000000") AFTER 510ns, 
 ("00000000000000000000000000000000") AFTER 520ns, 
 ("00000000000000000000000000000000") AFTER 530ns, 
 ("00000000000000000000000000000000") AFTER 540ns, 
 ("00000000000000000000000000000000") AFTER 550ns; 
 
 En_tb <= '1';
 RST_tb <= '1' , '0' AFTER 8ns;
 
 Process_3: Process(H_t_tb,C_t_tb)
    VARIABLE outline_C_t : LINE;
    VARIABLE outline_H_t : LINE;
    VARIABLE linenumber : INTEGER := 0;
    FILE C_t_file : TEXT OPEN write_mode IS "C:\Users\bpa4hi\LSTM\C_t.txt";
    FILE H_t_file : TEXT OPEN write_mode IS "C:\Users\bpa4hi\LSTM\H_t.txt";
    BEGIN 
            write(outline_C_t,TO_INTEGER(SIGNED(C_t_tb)));
            writeline(C_t_file, outline_C_t);
            write(outline_H_t,TO_INTEGER(SIGNED(H_t_tb)));
            writeline(H_t_file, outline_H_t);
    END PROCESS;
 END Behavioral;
