----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09/11/2017 01:30:01 PM
-- Design Name: 
-- Module Name: Tanh - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.ALL;
LIBRARY WORK;
USE WORK.Generic_size_of_matrices_pkg.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

ENTITY Sigmoid IS
       PORT ( Din: IN Fixed_Point;
              Dout: OUT Fixed_Point);
        
END Sigmoid;

ARCHITECTURE Behavioral OF Sigmoid IS

SIGNAL TEMP : SIGNED(31 DOWNTO 0);
BEGIN

TEMP <= SIGNED(Din);

 PROCESS(TEMP)
 BEGIN
  CASE (TO_INTEGER(TEMP)) IS   
          WHEN -2147483648 TO -262144 => Dout <= "00000000000000000000010010011011";
          WHEN -262143 TO -255590 => Dout <="00000000000000000000010100010101";
          WHEN -255589 TO -249036 => Dout <="00000000000000000000010110011011";
          WHEN -249035 TO -242483 => Dout <="00000000000000000000011000101110";
          WHEN -242482 TO -235929 => Dout <="00000000000000000000011011010000";
          WHEN -235928 TO -229376 => Dout <="00000000000000000000011110000010";
          WHEN -229375 TO -222822 => Dout <="00000000000000000000100001000101";
          WHEN -222821 TO -216268 => Dout <="00000000000000000000100100011100";
          WHEN -216267 TO -209715 => Dout <="00000000000000000000101000000111";
          WHEN -209714 TO -203161 => Dout <="00000000000000000000101100001010";
          WHEN -203160 TO -196608 => Dout <="00000000000000000000110000100101";
          WHEN -196607 TO -190054 => Dout <="00000000000000000000110101011010";
          WHEN -190053 TO -183500 => Dout <="00000000000000000000111010101101";
          WHEN -183499 TO -176947 => Dout <="00000000000000000001000000100000";
          WHEN -176946 TO -170393 => Dout <="00000000000000000001000110110100";
          WHEN -170392 TO -163840 => Dout <="00000000000000000001001101101100";
          WHEN -163839 TO -157286 => Dout <="00000000000000000001010101001011";
          WHEN -157285 TO -150732 => Dout <="00000000000000000001011101010100";
          WHEN -150731 TO -144179 => Dout <="00000000000000000001100110001010";
          WHEN -144178 TO -137625 => Dout <="00000000000000000001101111101110";
          WHEN -137624 TO -131072 => Dout <="00000000000000000001111010000101";
          WHEN -131071 TO -124518 => Dout <="00000000000000000010000101001111";
          WHEN -124517 TO -117964 => Dout <="00000000000000000010010001010001";
          WHEN -117963 TO -111411 => Dout <="00000000000000000010011110001100";
          WHEN -111410 TO -104857 => Dout <="00000000000000000010101100000001";
          WHEN -104856 TO -98304 => Dout <= "00000000000000000010111010110100";
          WHEN -98303 TO -91750 => Dout <= "00000000000000000011001010100101";
          WHEN -91749 TO -85196 => Dout <= "00000000000000000011011011010100";
          WHEN -85195 TO -78643 => Dout <= "00000000000000000011101101000010";
          WHEN -78642 TO -72089 => Dout <= "00000000000000000011111111101111";
          WHEN -72088 TO -65536 => Dout <= "00000000000000000100010011011010";
          WHEN -65535 TO -58982 => Dout <= "00000000000000000100101000000000";
          WHEN -58981 TO -52428 => Dout <= "00000000000000000100111101011110";
          WHEN -52421 TO -45875 => Dout <= "00000000000000000101010011110010";
          WHEN -45874 TO -39321 => Dout <="00000000000000000101101010110111";
          WHEN -39320 TO -32768 => Dout <= "00000000000000000110000010100111";
          WHEN -32767 TO -26214 => Dout <= "00000000000000000110011010111101";
          WHEN -26213 TO -19660 => Dout <= "00000000000000000110110011110010";
          WHEN -19659 TO -13107 => Dout <= "00000000000000000111001100111111";
          WHEN -13106 TO -6553 => Dout <="00000000000000000111100110011011";
          WHEN -6552 TO -1 => Dout <="00000000000000000111111110011011";
          WHEN   0 => Dout <=  "00000000000000001000000000000000"; --   A = 0
          WHEN 1 TO 6554 => Dout <="00000000000000001000011001100110";
          WHEN 6555 TO 13108 => Dout <="00000000000000001000110011000010";
          WHEN 13109 TO 19661 => Dout <= "00000000000000001001001100001111";
          WHEN 19662 TO 26215 => Dout <="00000000000000001001100101000100";
          WHEN 26216 TO 32768 => Dout <="00000000000000001001111101011010";
          WHEN 32769 TO 39322 => Dout <="00000000000000001010010101001010";
          WHEN 39323 TO 45876 => Dout <="00000000000000001010101100001111";
          WHEN 45877 TO 52429 => Dout <="00000000000000001011000010100011";
          WHEN 52430 TO 58983 => Dout <="00000000000000001011011000000001";
          WHEN 58984 TO 65536 => Dout <="00000000000000001011101100100111";
          WHEN 65537 TO 72090 => Dout <="00000000000000001100000000010010";
          WHEN 72091 TO 78644 => Dout <="00000000000000001100010010111111";
          WHEN 78645 TO 85197 => Dout <="00000000000000001100100100101101";
          WHEN 85198 TO 91751 => Dout <="00000000000000001100110101011100";
          WHEN 91752 TO 98304 => Dout <="00000000000000001101000101001101";
          WHEN 98305 TO 104858 => Dout <="00000000000000001101010100000000";
          WHEN 104859 TO 111412 => Dout <="00000000000000001101100001110101";
          WHEN 111413 TO 117965 => Dout <="00000000000000001101101110110000";
          WHEN 117966 TO 124519 => Dout <="00000000000000001101111010110010";
          WHEN 124520 TO 131072 => Dout <="00000000000000001110000101111100";
          WHEN 131073 TO 137626 => Dout <="00000000000000001110010000010011";
          WHEN 137627 TO 144180 => Dout <="00000000000000001110011001110111";
          WHEN 144181 TO 150733 => Dout <="00000000000000001110100010101101";
          WHEN 150734 TO 157287 => Dout <="00000000000000001110101010110110";
          WHEN 157288 TO 163840 => Dout <="00000000000000001110110010010101";
          WHEN 163841 TO 170394 => Dout <="00000000000000001110111001001101";
          WHEN 170395 TO 176948 => Dout <="00000000000000001110111111100001";
          WHEN 176949 TO 183501 => Dout <="00000000000000001111000101010100";
          WHEN 183502 TO 190055 => Dout <="00000000000000001111001010100111";
          WHEN 190056 TO 196608 => Dout <="00000000000000001111001111011100";
          WHEN 196609 TO 203162 => Dout <="00000000000000001111010011110111";
          WHEN 203163 TO 209716 => Dout <="00000000000000001111010111111010";
          WHEN 209717 TO 216269 => Dout <="00000000000000001111011011100101";
          WHEN 216270 TO 222823 => Dout <="00000000000000001111011110111100";
          WHEN 222824 TO 229376 => Dout <="00000000000000001111100001111111";
          WHEN 229377 TO 235930 => Dout <="00000000000000001111100100110001";
          WHEN 235931 TO 242484 => Dout <="00000000000000001111100111010011";
          WHEN 242485 TO 249037 => Dout <="00000000000000001111101001100110";
          WHEN 249038 TO 255591 => Dout <="00000000000000001111101011101100";
          WHEN 255592 TO 262144 => Dout <="00000000000000001111101101100110";
          WHEN OTHERS =>  Dout <=    "00000000000000001111101101100110"; 
      END CASE;
END PROCESS;

END Behavioral;
